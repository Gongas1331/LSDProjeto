library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity MaqLavar is
end MaqLavar;

architecture Shell of MaqLavar is
end Shell;